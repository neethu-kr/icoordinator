<?php
global $langArray;
$brand_name = getenv('BRAND_NAME');
$langArray = array(
    "files_not_uploaded" => "Filerna har inte laddats upp",
    "files_not_uploaded_msg" => "Dina filer som skickades med inkommande e-post har inte laddats upp. Vänligen kontakta portaladministratören för mer information.",
    "files_not_uploaded_email_msg" => "Dina filer som skickades med inkommande e-post har inte laddats upp. Kontrollera den e-postadress du skickat till",
    "files_uploaded" => "Filerna har laddats upp.",
    "files_uploaded_msg" => "Dina filer som skickades med inkommande e-post har laddats upp.",
    "files" => "Filer",
    "password_reset_success_msg" => "Ett nytt automatgenererat lösenord till ditt ".$brand_name."-konto har skapats.",
    "new_password" => "Nytt lösenord",
    "portal_invitation_greeting" => "Du har blivit inbjuden till ".$brand_name,
    "portal_invitation_msg" => "*|INVITED_BY_NAME|* har bjudit in dig att arbeta på följande portal",
    "accept_invitation" => "Acceptera inbjudan",
    "notification_report" => "Notifieringsrapport",
    "shared_file_notification_greeting" => "En fil har delats med dig",
    "shared_file_notification_msg" => "*|USER_NAME|* har delat följande fil med dig",
    "shared_files_notification_greeting" => "*|USER_NAME|* har delat mappinformation med dig",
    "shared_files_notification_msg" => "",
    "message" => "Meddelande",
    "shared_folder_notification_greeting" => "En mapp har delats med dig",
    "shared_folder_notification_msg" => "*|USER_NAME|* har delat följande mapp med dig",
    "sign_up_confirm_greeting" => "Verifiera ditt e-postmeddelande för att börja använda ". $brand_name,
    "welcome_to_brand" => "Välkommen till ".$brand_name,
    "sign_up_comfirm_msg" => "Verifiera din e-postadress för att komma igång. Vi gör detta som en säkerhetsåtgärd för att verifiera dina uppgifter",
    "verify_email" => "Verifiera e-post",
    "invitation_greeting" => "Du har blivit inbjuden till ".$brand_name,
    "invitation_msg" => "*|INVITED_BY_NAME|* har bjudit in dig till ".$brand_name." för att arbeta i följande portal",
    "invitation_accepted_msg" => "Du har nu accepterat inbjudan att arbeta i portalen ",
    "here_are_your_credentials" => "Här är dina uppgifter",
    "login" => "Logga in",
    "password" => "Lösenord",
    "start_collaborating_msg" => "Gå till *|WEB_BASE_URL|* för att logga in och börja samarbeta.",
    "thank_you_for_using_brand" => "Tack för att du använder ".$brand_name,
    "brand_account_created" => "Ditt ".$brand_name." konto skapades",
    "inbound_unexpected_server_error" => "Ingående epost: Oväntat serverfel",
    "inbound_successful_upload" => "Ingående epost: Filen laddades upp",
    "inbound_wrong_email" => "Ingående epost: Felaktig epostadress",
    "password_reset_success" => "Ett nytt automatgenererat lösenord har skapats",
    "invitation_to_portal" => "Inbjudan till portalen *|PORTAL_NAME|*",
    "brand_notification_report" => $brand_name . " prenumerationsrapport",
    "notification_file_was_shared" => "Filen *|FILE_NAME|* har delats med dig",
    "notification_files_were_shared" => "Filer från *|WORKSPACE_NAME|* i mappen *|FOLDER_NAME|* delades med dig",
    "notification_folder_was_shared" => "Mappen *|FOLDER_NAME|* har delats med dig",
    "complete_brand_signup" => "Vänligen slutför registreringen av ditt " . $brand_name . "-konto",
    "invitation_to_brand" => "Inbjudan till " . $brand_name,
    "file_created_by" => "Filen skapades av",
    "file_updated_by" => "Filen uppdaterades av",
    "file_deleted_by" => "Filen togs bort av",
    "file_uploaded_by" => "Filen laddades upp av",
    "file_new_version_uploaded_by" => "Ny version laddades upp av",
    "portal" => "Portal",
    "workspace" => "Arbetsyta",
    "new_workspace" => "Ny arbetsyta",
    "copy_workspace_subject" => "Kopiera arbetsyta: Arbetsytan skapades",
    "copy_workspace_header" => "Arbetsytan skapades",
    "copy_workspace_workspace_created" => "Arbetsytan skapad via kopiera arbetsyta-funktionaliteten är nu redo att användas."
);